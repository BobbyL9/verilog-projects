module regfile
(
    input logic clk, we3,
    input logic [4:0] a1, a2, a3,
    input logic wd3,
    output logic rd1,
    output logic rd2
);

//regfile rf(clk, regwrite, instr[19:15], instr[24:20], instr[11:7], result, srca, writedata);


endmodule
